/*
 * GPU_GEO_tb.sv, for ModelSim and ***NEW Active-HDL.
 *
 * Features control from a source ASCII text file script,
 * and a 256 color .BMP picture file generator.
 * Tested on free Altera ModelSim 10 & 20.  Built in parameter
 * (USE_ALTERA_IP) when disabled prevents the use of any Altera specific IP functions.
 *
 * Written by Brian Guralnick.
 *
 * v 0.6.001   Feb 01, 2021
 *
 * To setup simulation, Start Modelsim, Then go to 'File - Change Directory' and select this files directory. 
 * Then in the transcript, type:
 * do setup_ms.do
 * (or if you want to enable the Altera megafunction IP, LPM_MULT & SCFIFO)
 * do setup_altera.do
 * 
 * To change the 'TB_COMMAND_SCRIPT_FILE' source script file string and re-run the simulation, type:
 *
 * do test_8bitfont.do
 * do test_45deg.do
 * do test_art.do
 * do test_blitter.do
 * do test_blitter_hires.do
 * do test_vwait.do
 *
 *
 *****************************************************************************
 * For Active-HDL (Comes with Lattice Diamond FPGA development environment.)
 *****************************************************************************
 *
 * Go to 'File - New / Design'
 *        Create an empty design.
 *        Choose Verilog for HDL language, ignore 'Target Technology'.
 *        Type in 'GPU_GEO_tb' for design name.
 *        Next/Finish.
 *        
 * Unzip all the files directly into the 'src' directory inside the 'GPU_GEO_tb' folder.
 * In the console, type:
 *
 * do setup_active-hdl.do
 *
 * *** The result 'xxxx.bmp' and 'GEO_tb_command_results.txt' files generated by
 *     the simulation will be located in the main 'GPU_GEO_tb' folder.
 *
 * Active-HDL does not support the changing of a string in a .sv file,
 * so to run the different tb ASCII script demos, you need to copy the:
 *
 * GEO_tb_art.txt
 * GEO_tb_Blitter.txt
 * GEO_tb_Blitter_hires.txt
 * GEO_tb_45deg_zilog.txt
 * GEO_tb_8bit_font.txt
 * GEO_tb_vwait.txt
 *
 * over the 'GEO_tb_command_list.txt' file, then do a restart & run simulation.
 *
 */

`timescale 1 ns/ 1 ns // 1 ns steps, 1 ns precision.

module GPU_GEO_tb 
#(
parameter int BITS_RES                  = 12,
parameter bit USE_ALTERA_IP             = 0,
parameter int PIXIE_MEM_ADR             = 20
)();
string TB_COMMAND_SCRIPT_FILE = "GEO_tb_command_list.txt";	 // Choose one of the following strings...
//string TB_COMMAND_SCRIPT_FILE = "GEO_tb_art.txt";
//string TB_COMMAND_SCRIPT_FILE = "GEO_tb_Blitter.txt";
//string TB_COMMAND_SCRIPT_FILE = "GEO_tb_Blitter_hires.txt";
//string TB_COMMAND_SCRIPT_FILE = "GEO_tb_45deg_zilog.txt";
//string TB_COMMAND_SCRIPT_FILE = "GEO_tb_8bit_font.txt";
//string TB_COMMAND_SCRIPT_FILE = "GEO_tb_vwait.txt";

// GPU_GEO_tb master controls
logic                     hse,vse;                 // Dummy Syncs for the V-wait command
logic                     clk,reset;
logic                     TB_cmd_ena;              // Strobe high to send the command to DUT_GEOFF.
logic [15:0]              TB_cmd_in;               // Contains the 16bit command

// DUT_GEOFF results
logic                     GEOFF_busy;              // Only send TB_cmd_ena when this status flag is low.
logic                     GEOFF_draw_cmd_rdy;
logic [35:0]              GEOFF_draw_cmd;

logic                     PAGET_cmd_rdy;
logic [39:0]              PAGET_cmd;

logic                     PIXIE_busy;
logic                     PIXIE_rd_req_a,PIXIE_rd_req_b,PIXIE_wr_ena;
logic [PIXIE_MEM_ADR-1:0] PIXIE_ram_addr;
logic [15:0]              PIXIE_ram_wr_data;
logic                     RAM_ctl_busy;                       // Tells PIXIE that the ram controller isn't ready to receive a command.
logic                     RAM_data_rdy_a,RAM_data_rdy_b;      // ram block read-request return
logic [15:0]              RAM_data_read;                      // ram block read data from 

logic                     PIXIE_col_rd_rst,PIXIE_col_wr_rst;  // PIXIE read/write collision detect reset
logic [7:0]               PIXIE_col_rd,PIXIE_col_wr ;

string                Script_CMD  = "" ; // Message line in waveform
logic [12:0]          Script_LINE = 0  ; // Message line in waveform
logic                 ENA_PIXIE   = 0  ;

logic unsigned [23:0] PAGER_base_adr[0:1]   = '{0,0}; // srce/dest base address.
logic unsigned [23:0] PAGER_base_width[0:1] = '{0,0}; // srce/dest bitmap width.
logic unsigned [ 7:0] PAGER_base_depth[0:1] = '{0,0}; // srce/dest bitmap depth.

wire unsigned [3:0]  GEOFF_cmd_cmd   = GEOFF_draw_cmd[35:32];
wire unsigned [7:0]  GEOFF_cmd_color = GEOFF_draw_cmd[31:24];
wire unsigned [11:0] GEOFF_cmd_y     = GEOFF_draw_cmd[23:12];
wire unsigned [11:0] GEOFF_cmd_x     = GEOFF_draw_cmd[11:0 ];
localparam bit [3:0] CMD_DRAW = 1;


wire unsigned [3:0]  PAGET_cmd_cmd   = PAGET_cmd[39:36];
wire unsigned [7:0]  PAGET_cmd_color = PAGET_cmd[35:28];
wire unsigned [3:0]  PAGET_cmd_depth = PAGET_cmd[27:24];
wire unsigned [3:0]  PAGET_cmd_bit   = PAGET_cmd[23:20];
wire unsigned [19:0] PAGET_cmd_addr  = PAGET_cmd[19:0 ];

logic GEOFF_busy_internal;

localparam CLK_MHz  = 100 ;
localparam period  = 1000/CLK_MHz ;    // Calculate the clk toggle rate.

localparam HS_PIXEL = 64 ;             // Make a dummy hsync pulse every 16 pixels.
localparam VS_PIXEL = 48 ;             // Make a dummy vsync pulse every 8  hsyncs.

integer h_cnt,v_cnt;

geometry_xy_plotter #(.USE_ALTERA_IP(USE_ALTERA_IP)) DUT_GEOFF (

   // inputs
   .clk            ( clk             ),
   .reset          ( reset           ),
   .fifo_cmd_ready ( TB_cmd_ena      ),
   .fifo_cmd_in    ( TB_cmd_in       ),
   .draw_busy      ( PIXIE_busy      ),
   .hse            ( hse             ),
   .vse            ( vse             ),

   //outputs
   .load_cmd       (                     ),        // HIGH when ready to receive next cmd_data[15:0] input
   .draw_cmd_rdy   ( GEOFF_draw_cmd_rdy  ),
   .draw_cmd       ( GEOFF_draw_cmd      ),
   .fifo_cmd_busy  ( GEOFF_busy          ),
   .processing     ( GEOFF_busy_internal ) );




pixel_address_generator #(.USE_ALTERA_IP(USE_ALTERA_IP)) DUT_PAGET (

    // inputs
    .clk           ( clk                 ),
    .reset         ( reset               ),
    .draw_cmd_rdy  ( GEOFF_draw_cmd_rdy  ),  // use _r, or _r2 to add a D-Clocked buffer between this section and the plotter.
    .draw_cmd      ( GEOFF_draw_cmd      ),  // use _r, or _r2 to add a D-Clocked buffer between this section and the plotter.
    .draw_busy     ( PIXIE_busy          ),

    // outputs
    .pixel_cmd_rdy ( PAGET_cmd_rdy       ),
    .pixel_cmd     ( PAGET_cmd           ) );



geo_pixel_writer DUT_PIXIE (

    // inputs
    .clk              ( clk              ),
    .reset            ( reset            ),
    .cmd_rdy          ( PAGET_cmd_rdy && ENA_PIXIE && !PIXIE_busy ),
    .cmd_in           ( PAGET_cmd        ),
    .rd_data_in       ( RAM_data_read    ),
    .rd_data_rdy_a    ( RAM_data_rdy_a   ),
    .rd_data_rdy_b    ( RAM_data_rdy_b   ),
    .ram_mux_busy     ( RAM_ctl_busy     ),
    .collision_rd_rst ( PIXIE_col_rd_rst ),
    .collision_wr_rst ( PIXIE_col_wr_rst ),

    // outputs
    .draw_busy        ( PIXIE_busy       ),
    .rd_req_a         ( PIXIE_rd_req_a   ),
    .rd_req_b         ( PIXIE_rd_req_b   ),
    .wr_ena           ( PIXIE_wr_ena     ),
    .ram_addr         ( PIXIE_ram_addr   ),
    .ram_wr_data      ( PIXIE_ram_wr_data),
    .collision_rd     ( PIXIE_col_rd     ),
    .collision_wr     ( PIXIE_col_wr     ),
    .PX_COPY_COLOUR   (                  ) );





// ***********************************************************************************************************
// ***********************************************************************************************************
// Setup global bitmap size and logic memory array.
//
localparam BMP_WIDTH  = 1024;
localparam BMP_HEIGHT = 1024;
logic [7:0] bitmap [0:BMP_WIDTH-1][0:BMP_HEIGHT-1];
logic       BW_BMP = 0;     // set to 1 for 256 shades of grey BMP.
//
// ***********************************************************************************************************
// ***********************************************************************************************************

// ***********************************************************************************************************
// ***********************************************************************************************************
// Setup emulated Altera lpm_ram block ram memory array 
//
logic [15:0]                GPU_RAM [0:((2**(PIXIE_MEM_ADR-1))-1)] = '{(2**(PIXIE_MEM_ADR-1)){0}}; // This is all the ram.
logic [(PIXIE_MEM_ADR-1):0] GPU_RAM_adr_in   = 0;
logic [(PIXIE_MEM_ADR-1):0] GPU_RAM_adr_rd   = 0;
logic [(PIXIE_MEM_ADR-1):0] GPU_RAM_data_in  = 0;
logic                       GPU_RAM_we       = 0;
logic                       gpu_ram_rdreq_a  = 0;
logic                       gpu_ram_rdreq_b  = 0;
logic                       gpu_ram_rdreq_ma = 0;
logic                       gpu_ram_rdreq_mb = 0;
//
// ***********************************************************************************************************
// ***********************************************************************************************************


logic       [7:0] WDT_COUNTER;          // Wait for 15 clocks or inactivity before forcing a simulation stop.
logic             WAIT_IDLE = 0;        // When high, insert a idle wait before every command.
localparam int    WDT_RESET_TIME = 24;  // Set tyhe WDT timeout clock cycles.
localparam int    SYS_IDLE_TIME = WDT_RESET_TIME-12; // Consider system idle after 12 clocks of inactivity.

// This logic creates 1 flag which goes high if any modules are doing anything, or they are busy.
// It is used for the watchdog timer and waiting for all operations to finish before doing things like save a .BMP image.
logic         busy_system ;
always_comb   busy_system = ( reset || TB_cmd_ena || GEOFF_busy || GEOFF_busy_internal || GEOFF_draw_cmd_rdy || PAGET_cmd_rdy || PIXIE_busy || PIXIE_rd_req_a || PIXIE_rd_req_b || PIXIE_wr_ena ) ;


initial 
begin 
clk              = 1'b1;
reset            = 1'b1;  // apply reset
WDT_COUNTER      = WDT_RESET_TIME  ; // Set the initial inactivity timer to maximum so that the code later-on wont immediately stop the simulation.
TB_cmd_ena       = 0;
TB_cmd_in        = 0;
hse              = 0;
vse              = 0;
h_cnt            = 0;
v_cnt            = 0;
RAM_ctl_busy     = 0;
RAM_data_rdy_a   = 0;
RAM_data_rdy_b   = 0;
RAM_data_read    = 0;
PIXIE_col_rd_rst = 0;
PIXIE_col_wr_rst = 0;
GPU_RAM [0:((2**(PIXIE_MEM_ADR-1))-1)] = '{(2**(PIXIE_MEM_ADR-1)){0}}; // This is all the ram.
GPU_RAM_adr_in   = 0;
GPU_RAM_adr_rd   = 0;
GPU_RAM_data_in  = 0;
GPU_RAM_we       = 0;
gpu_ram_rdreq_a  = 0;
gpu_ram_rdreq_b  = 0;
gpu_ram_rdreq_ma = 0;
gpu_ram_rdreq_mb = 0;
Script_CMD       = "";
Script_LINE      = 0;
ENA_PIXIE        = 0;

PAGER_base_adr[0:1]   = '{0,0}; // srce/dest base address.
PAGER_base_width[0:1] = '{0,0}; // srce/dest bitmap width.
PAGER_base_depth[0:1] = '{0,0}; // srce/dest bitmap depth.


#(period*2);
reset = 1'b0; // clear reset
#(period*2);

@(negedge clk); // Align to the negedge clock.
WDT_COUNTER = WDT_RESET_TIME;
execute_ascii_file(TB_COMMAND_SCRIPT_FILE); // Run the ASCII test bench script.

end 

// Always cycle clk logic at the period speed.
always #(period/2) clk = !clk;

// Create a watchdog inactivity countdown timer called running.
// When logic is busy or set to run, reset the timer to 16, otherwise
// decrement every clk cycle.
always @(posedge clk) WDT_COUNTER = (busy_system) ? WDT_RESET_TIME : (WDT_COUNTER-1'b1) ;   // Setup a simulation inactivity watchdog countdown timer.
always @(posedge clk) if (WDT_COUNTER==0) $stop;                             // Automatically stop the simulation if the inactivity timer reaches 0.


// Trap and plot GEOFF pixel write commands into bitmap buffer
always @(negedge clk) if (GEOFF_cmd_x>=0 && GEOFF_cmd_y>=0 && GEOFF_cmd_x<BMP_WIDTH && GEOFF_cmd_y<BMP_HEIGHT && (GEOFF_cmd_cmd==CMD_DRAW)) bitmap[GEOFF_cmd_x][GEOFF_cmd_y] = GEOFF_cmd_color;


// ***********************************************************************************************************
//Generate a dummy hse and vse sync pulses to test the vwait command.
// ***********************************************************************************************************
always @(negedge clk) begin
	hse = (h_cnt==0);
        vse = (v_cnt==0);
	if (h_cnt>=HS_PIXEL-1) begin
                      h_cnt = 0;
	              if (v_cnt>=VS_PIXEL-1) v_cnt = 0;
                      else v_cnt++;
        end else h_cnt++;
end
// ***********************************************************************************************************
// Emulate Altera lpm_ram block ram memory array with 1 clock write, 2 clock read, dont care read while write result
// ***********************************************************************************************************
always @(posedge clk) begin

// latch command from PIXIE
GPU_RAM_adr_in  <= PIXIE_ram_addr;
GPU_RAM_we      <= PIXIE_wr_ena;
GPU_RAM_data_in <= PIXIE_ram_wr_data;
gpu_ram_rdreq_a <= PIXIE_rd_req_a;
gpu_ram_rdreq_b <= PIXIE_rd_req_b;

// Write data...
if (GPU_RAM_we) GPU_RAM[(GPU_RAM_adr_in>>1)] <= GPU_RAM_data_in ;

// Read data 1 additional clock later
GPU_RAM_adr_rd   <= GPU_RAM_adr_in;
gpu_ram_rdreq_ma <= gpu_ram_rdreq_a;
gpu_ram_rdreq_mb <= gpu_ram_rdreq_b;

// Send read result back to PIXIE
RAM_data_read    <= GPU_RAM[(GPU_RAM_adr_rd>>1)];
RAM_data_rdy_a   <= gpu_ram_rdreq_ma;
RAM_data_rdy_b   <= gpu_ram_rdreq_mb;

end
// ***********************************************************************************************************



// ***********************************************************************************************************
// ***********************************************************************************************************
// ***********************************************************************************************************
//
// End of test-bench.
//
// Next, 'task' programs:
//
// save_bmp_256( "bmp_file_name.bmp" , <bw_nocolor> );      // saves a 256 color BMP picture.
// execute_ascii_file("<source file name">);                // Executes the command ASCII file, decodes the '@' command string
//
// draw_ellipse(*src, *dest, fill, first quad, end quad);     // reads source file for coordinates, then runs the ellipse generator
// clear_bitmap(integer xs, integer ys, byte unsigned color); // clears the logic array bitmap to byte 'color'
// task send_rst();                                           // pulses the reset line.
//
// ***********************************************************************************************************
// ***********************************************************************************************************
// ***********************************************************************************************************





// ***********************************************************************************************************
// ***********************************************************************************************************
// ***********************************************************************************************************
// Simple 256 color BMP save algorithm.
// To call task:
//
// save_bmp_256( "bmp_file_name.bmp" , <bw_nocolor>, <xsize>, <ysize>, use_pixie, pixie_dest );
//
// If (bw_nocolor=1), the result bitmap will be 256 shades of grey from 0=black to 255=white.
// If (bw_nocolor=0), the result bitmap will have a dummy color palette.
//
// 
// logic array 'bitmap' must be declared at the top of the test-bench module like this:
// logic   [7:0] bitmap [0:BMP_WIDTH-1][0:BMP_HEIGHT-1];
//
// When rendering into the array 'bitmap', it is recommended you use range checks such as:
//
// if (X_coord>=0 && Y_coord>=0 && X_coord<BMP_WIDTH && Y_coord<BMP_HEIGHT) bitmap[X_coord][Y_coord] = draw_color;
// 
// ***********************************************************************************************************
//  BMP Header
// 16 bit string "BM", first 2 bytes in file, but ignored everywhere else...
// 32 bit, offset 0002, Full size of BMP file in bytes. = 54(header not including 'BM') + 1024(palette) + (BMP_WIDTH(word padded)*BMP_HEIGHT)
// 32 bit, offset 0006, Dummy 32'h0000
// 32 bit, offset 000A, First byte of where the the bitmap data begins. - 1078 = 54(header)+1024(palette)
// 32 bit, offset 000E, Size of header in bytes.   Must be 40
// 32 bit, offset 0012, BMP_WIDTH
// 32 bit, offset 0016, BMP_HEIGHT
// 16 bit, offset 001A, Number of color planes. Must be     1
// 16 bit, offset 001C, Color depth. Must be 1,4,8,16,24,32 8 = 8 bit per pixel
// 32 bit, offset 001E, Compression method used.            0 = none.
// 32 bit, offset 0022, Image size in bytes.                  = BMP_row_size*BMP_HEIGHT   (Remember 4 byte per line padding) 
// 32 bit, offset 0026, Horizontal res, pixel/meter,     2835 = 72 pixels per inch
// 32 bit, offset 002A, Vertical   res, pixel/meter,     2835 = 72 pixels per inch
// 32 bit, offset 002E, Number of colors in palette.     256.
// 32 bit, offset 0032, Number of important colors used. 256.
// ***********************************************************************************************************
// ***********************************************************************************************************

task save_bmp_256(string bmp_file_name,bit bw_nocolor,integer width, integer height, bit use_pixie, bit pd);
begin

    integer unsigned        fout_bmp_pointer, BMP_file_size,BMP_row_size,r;
    logic   unsigned [31:0] BMP_header[0:12];

                            BMP_row_size  = 32'(width) & 32'hFFFC; // When saving a bitmap, the row size/width must be
if ((width & 32'd3) !=0)    BMP_row_size  = BMP_row_size + 4;      // padded to chunks of 4 bytes.

    fout_bmp_pointer= $fopen(bmp_file_name,"wb");
    if (fout_bmp_pointer==0)
    begin
       $display("Could not open file '%s' for writing",bmp_file_name);
       $stop;     
    end
    $display(" *************************************************************** ");
    $display(" ****** Saving bitmap '%s'. ********** ",bmp_file_name);
    $display(" *************************************************************** ");


BMP_file_size    = (54+1024+(BMP_row_size*height));

BMP_header[0:12] = '{BMP_file_size,0,1078,40,width,height,{16'd8,16'd1},0,(BMP_row_size*height),2835,2835,256,256};

//$fwrite(fout_bmp_pointer,"BM%u",BMP_header); //  Not compatible with Lattice Active_HDL.
$fwrite(fout_bmp_pointer,"BM");
for (int i =0 ; i <13 ; i++ ) $fwrite(fout_bmp_pointer,"%u",BMP_header[i]); // Better compatibility with Lattice Active_HDL.


    //  Save 256 color .bmp palette
    if (!bw_nocolor) for (int i=0 ; i<256 ; i++)  $fwrite(fout_bmp_pointer,"%c%c%c%c",8'({i[3:0],i[3:0]}),8'({i[5:2],i[5:2]}),8'({i[7:4],i[7:4]}),8'h00);// Generate a dummy colorized palette
    // This makes the palette go from color 0=black to 255=100% white.
    else             for (int i=0 ; i<256 ; i++)  $fwrite(fout_bmp_pointer,"%u",({8'h00,8'(i),8'(i),8'(i)})); // Generate a monochrome 256 shade grey palette

    //  Save BMP_WIDTHxBMP_HEIGHT .bmp image.
    for (int y=height-1;y>=0;y--) begin
                                  for (int x=0;x<width;x+=4) begin
                                                             // Save GEOFF XY plotter pixel output
                                                             if (!use_pixie) $fwrite(fout_bmp_pointer,"%u",{bitmap[x+3][y],        bitmap[x+2][y],        bitmap[x+1][y],        bitmap[x][y]}) ;
                                                             // Save GPU ram image output
                                                             else            $fwrite(fout_bmp_pointer,"%u",{pixie_pixel(pd,x+3,y), pixie_pixel(pd,x+2,y), pixie_pixel(pd,x+1,y), pixie_pixel(pd,x,y)}) ;
                                                             end
                                  end


    $fclose(fout_bmp_pointer);
end

endtask


// ***********************************************************************************************************
// ***********************************************************************************************************
// ***********************************************************************************************************
// task execute_ascii_file(<"source ASCII file name">);
// 
// Opens the ASCII file and scans for the '@' symbol.
// After each '@' symbol, a string is read as a command function.
// Each function then goes through a 'case(command_in)' which then executes the appropriate function.
//
// ***********************************************************************************************************
// ***********************************************************************************************************
// ***********************************************************************************************************

task execute_ascii_file(string source_file_name);
 begin
    integer unsigned fin_pointer,fout_pointer,fin_running,r,x,y,z;
    string  command_in,message_string,destination_file_name,bmp_file_name,msg;

    byte    unsigned    char        ;
    byte    unsigned    draw_color  ;
    integer unsigned    line_number ;

    line_number  = 1;
    fout_pointer = 0;
    fin_pointer  = 0;

    fin_pointer= $fopen(source_file_name, "r");
    if (fin_pointer==0)
    begin
       $display("Could not open file '%s' for reading",source_file_name);
       $stop;     
    end

while (fin_pointer!=0 && ! $feof(fin_pointer)) begin // Continue processing until the end of the source file.

  char = 0;
  while (char != "@" && ! $feof(fin_pointer) && fin_pointer!=0 ) begin // scan for the @ character until end of source file.
  char = $fgetc(fin_pointer);
  if (char==0 || fin_pointer==0 )  $stop;                               // something went wrong
  if (char==10) line_number = line_number + 1;       // increment the internal source file line counter.
  end


if (! $feof(fin_pointer) && fin_pointer!=0) begin  // if not end of source file retrieve command string

  r = $fscanf(fin_pointer,"%s",command_in); // Read in the command string after the @ character.
  if (fout_pointer!=0) $fwrite(fout_pointer,"Line#%d, ",13'(line_number)); // :pg the executed command line number.

  case (command_in) // select command string.

  "SET_XY"      : script_set_xy(fin_pointer,fout_pointer,line_number);

  "SET_MAX_XY"  : max_xy(fin_pointer,fout_pointer,line_number);

  "SET_PAGET"   : set_paget(fin_pointer,fout_pointer,line_number);

  "DRAW"        : draw(fin_pointer,fout_pointer,line_number);       // draws the selected shape.

  "BLIT"        : blit(fin_pointer,fout_pointer,line_number);       // Executes blitter functions.

  "VWAIT"       : vwait(fin_pointer,fout_pointer,line_number);      // Executes the wait interrupt function.

  "SEND_CMD"    : begin
                 r = $fscanf(fin_pointer,"%h",z);
                 send_cmd(z,"SEND_CMD",line_number,fout_pointer);          // sends the command to the DUT_GEOFF
                 if (fout_pointer!=0) $fwrite(fout_pointer,"Sending command %h.\n",16'(z));
                 end

  "ENA_PIXIE"    : begin
                 r = $fscanf(fin_pointer,"%d",ENA_PIXIE);
                 cmd_null( (ENA_PIXIE ? "PIXIE Enabled. ":"Pixie Disabled.") );    // sends dummy text to the waveform display
                 cmd_null( (ENA_PIXIE ? "PIXIE Enabled. ":"Pixie Disabled.") );    // sends dummy text to the waveform display
                 if (fout_pointer!=0) $fwrite(fout_pointer,"%s.\n",(ENA_PIXIE ? "PIXIE Enabled. ":"Pixie Disabled."));
                 end

  "WAIT_IDLE"    : begin
                 r = $fscanf(fin_pointer,"%d",WAIT_IDLE);
                 cmd_null( (WAIT_IDLE ? "Wait Idle ON. ":"Wait Idle OFF.") );    // sends dummy text to the waveform display
                 cmd_null( (WAIT_IDLE ? "Wait Idle ON. ":"Wait Idle OFF.") );    // sends dummy text to the waveform display
                 if (fout_pointer!=0) $fwrite(fout_pointer,"%s.\n",(WAIT_IDLE ? "Wait Idle ON. ":"Wait Idle OFF."));
                 end

  "RESET"      : begin
                 send_rst("RESET",line_number);                                          // pulses the reset signal for 1 clock.
                 if (fout_pointer!=0) $fwrite(fout_pointer,"Sending a reset to the entire system.\n");
                 end

  "LOAD_GPU_RAM" : load_gpu_ram(fin_pointer,fout_pointer,line_number,0);
  "SAVE_GPU_RAM" : save_gpu_ram(fin_pointer,fout_pointer,line_number,0);


  "CLR_GPU_RAM" : begin
                 wait_idle();
                 GPU_RAM [0:((2**(PIXIE_MEM_ADR-1))-1)] = '{(2**(PIXIE_MEM_ADR-1)){0}}; // This is all the ram.

                 $sformat(message_string,"Clear CLR_GPU_RAM.",draw_color);
                 cmd_null(message_string);
                 cmd_null(message_string);
                 if (fout_pointer!=0) $fwrite(fout_pointer,"%s\n",message_string);
                 end

  "CLR_BMP"    : begin
                 wait_idle();
                 r = $fscanf(fin_pointer,"%d",draw_color);
                 clear_bitmap(BMP_WIDTH,BMP_HEIGHT,draw_color);       // clears the 'bitmap' to a fixed color.

                 $sformat(message_string,"Clear GEOFF bitmap to color %d.",draw_color);
                 cmd_null(message_string);
                 cmd_null(message_string);
                 if (fout_pointer!=0) $fwrite(fout_pointer,"%s\n",message_string);
                 end

  "SAVE_GEO_BMP" : begin

                 wait_idle();

                 r = $fscanf(fin_pointer,"%s%d%d%d",bmp_file_name,x,y,BW_BMP); 
                   if (destination_file_name != "") begin
                       Script_LINE = line_number;
                       $sformat(message_string,"Save_GEO_BMP (%d,%d), %s",12'(x),12'(y),(BW_BMP ? "B&W.  ":"Color."));
                       cmd_null(message_string);
                       cmd_null(message_string);
                       if (fout_pointer!=0) $fwrite(fout_pointer,"%s\n",message_string);
                       save_bmp_256(bmp_file_name,BW_BMP,x,y,0,0);                                                            // Save the BMP image.
                   end else begin
                    $sformat(message_string,"\nInvalid file name for SAVE_GEO_BMP command.\n");
                    $display("%s",message_string);
                    $fclose(fin_pointer);
                    if (fout_pointer!=0) $fwrite(fout_pointer,"%s",message_string);
                    if (fout_pointer!=0) $fclose(fout_pointer);
                    $stop;
                   end
                 end

  "SAVE_PIXIE_BMP" : begin

                 wait_idle();

                 r = $fscanf(fin_pointer,"%s%s%d%d%d",bmp_file_name,msg,x,y,BW_BMP);
                       z=0;
                       if (msg[0]=="d" || msg[0]=="D") z=1;
 
                   if (destination_file_name != "") begin
                       Script_LINE = line_number;
                       $sformat(message_string,"Save_PIXIE_BMP %s (%d,%d), %s",(z ? "dest":"src "),13'(x),13'(y),(BW_BMP ? "B&W.  ":"Color."));
                       cmd_null(message_string);
                       if (fout_pointer!=0) $fwrite(fout_pointer,"%s\n",message_string);
                       save_bmp_256(bmp_file_name,BW_BMP,x,y,1,z);                                                            // Save the BMP image.
                   end else begin
                    $sformat(message_string,"\nInvalid file name for SAVE_PIXIE_BMP command.\n");
                    $display("%s",message_string);
                    $fclose(fin_pointer);
                    if (fout_pointer!=0) $fwrite(fout_pointer,"%s",message_string);
                    if (fout_pointer!=0) $fclose(fout_pointer);
                    $stop;
                   end
                 end

  "LOG_FILE"   : begin                                                  // begin logging the results.
                   if (fout_pointer==0) begin
                   r = $fscanf(fin_pointer,"%s",destination_file_name); // Read file name for the log file
                     fout_pointer= $fopen(destination_file_name,"w");   // Open that file name for writing.
                     if (fout_pointer==0) begin
                          $display("\nCould not open log file '%s' for writing.\n",destination_file_name);
                          $stop;
                     end else begin
                     $fwrite(fout_pointer,"Log file requested in '%s' at line#%d.\n\n",source_file_name,13'(line_number));
                     end
                   end else begin
                     $sformat(message_string,"\n*** Error in command script at line #%d.\n    You cannot open a LOG_FILE since the current log file '%s' is already running.\n    You must first '@END_LOG_FILE' if you wish to open a new log file.\n",13'(line_number),destination_file_name);
                     $display("%s",message_string);
                     $fclose(fin_pointer);
                     if (fout_pointer!=0) $fwrite(fout_pointer,"%s",message_string);
                     if (fout_pointer!=0) $fclose(fout_pointer);
                     $stop;
                   end
                 end

  "END_LOG_FILE" : if (fout_pointer!=0)begin                           // Stop logging the commands and close the current log file.
                       $sformat(message_string,"@%s command at line number %d.\n",command_in,13'(line_number));
                       $display("%s",message_string);
                       $fwrite(fout_pointer,"%s",message_string);
                       $fclose(fout_pointer);
                       fout_pointer = 0;
                   end

  "STOP"       :  begin // force a temporary stop.
                  $sformat(message_string,"@%s command at line number %d.\nType 'Run -All' to continue.",command_in,13'(line_number));
                  $display("%s",message_string);
                  if (fout_pointer!=0) $fwrite(fout_pointer,"%s",message_string);
                  $stop;
                  end

  "END"        :  begin // force seek to the end of the source file.

                 wait_idle();

                  $sformat(message_string,"@%s command at line number %d.\n",command_in,13'(line_number));
                  $display("%s",message_string);
                  $fclose(fin_pointer);
                  if (fout_pointer!=0) $fwrite(fout_pointer,"%s",message_string);
                  fin_pointer = 0;
                  end

  default      :  begin // Unknown command
                  $sformat(message_string,"Source ASCII file '%s' has an unknown command '@%s' at line number %d.\nProcessign stopped due to error.\n",source_file_name,command_in,13'(line_number));
                  $display("%s",message_string);
                  if (fout_pointer!=0) $fwrite(fout_pointer,"%s",message_string);
                  $stop;
                  end
  endcase

end // if !end of source file

end// while not eof


// Finished reading source file.  Close files and stop.
wait_idle();
$sformat(message_string,"\nEnd of command source ASCII file '%s'.\n%d lines processed.\n",source_file_name,13'(line_number));
$display("%s",message_string);
$fclose(fin_pointer);
if (fout_pointer!=0) $fwrite(fout_pointer,"%s",message_string);
if (fout_pointer!=0) $fclose(fout_pointer);
end
endtask







// ***********************************************************************************************************
// ***********************************************************************************************************
// ***********************************************************************************************************
// task clear_bitmap (integer xs, integer ys, byte unsigned color);
// 
// Clears the bitmap logic array with the 'color'
//
// ***********************************************************************************************************
// ***********************************************************************************************************
// ***********************************************************************************************************

task clear_bitmap (integer xs, integer ys, byte unsigned color);
begin

for(int y=0;y<ys;y++) begin
                      for(int x=0;x<xs;x++) bitmap [x][y]=color; 
                      end
end
endtask

// ***********************************************************************************************************
// task send_rst();
// sends a reset.
// ***********************************************************************************************************
task send_rst(string msg, integer ln);
begin
  if (msg != "") Script_CMD  = msg;
  if (msg != "") Script_LINE = ln;
reset = 1;
@(negedge clk); 
reset = 0;
@(negedge clk); 
//cmd_null( "" ); // Waits a clock & Leaves a clear space on the waveform
WDT_COUNTER = WDT_RESET_TIME;
end
endtask

// ***********************************************************************************************************
// task cmd_null( string  msg );
// Clears commands and inserts a script text
// ***********************************************************************************************************
task cmd_null( string msg );
begin
  wait_geoff(); // wait for busy to clear
  Script_CMD  = msg;
  @(negedge clk);
WDT_COUNTER = WDT_RESET_TIME;
end
endtask
// ***********************************************************************************************************
// task wait_geoff();
// Wait for DUT_GEOFF input buffer ready.
// ***********************************************************************************************************
task wait_geoff();
begin
  while (GEOFF_busy) @(negedge clk); // wait for busy to clear
end
endtask
// ***********************************************************************************************************
// task wait_idle();
// Wait for DUT_GEOFF the entire geometry system to become idle.
// needed before saving bitmaps or to space out commands.
// ***********************************************************************************************************
task wait_idle();
begin
Script_CMD = "Wait for all drawing to finish.";
  while (WDT_COUNTER > SYS_IDLE_TIME) @(negedge clk); // wait for busy to clear
  WDT_COUNTER          = WDT_RESET_TIME ; // Reset the watchdog timer.
end
endtask
// ***********************************************************************************************************
// task send_cmd( int cmd );
// sends a command.
// ***********************************************************************************************************
task send_cmd( int cmd, string msg, integer ln, integer dest );
begin
  logic unsigned [7:0] bh,bl;
  bh = cmd[15:8];
  bl = cmd[7:0];
  wait_geoff(); // wait for busy to clear
  TB_cmd_ena = 1;
  TB_cmd_in  = 16'(cmd);
  if (msg != "") Script_CMD  = msg;
  if (msg != "") Script_LINE = ln;
  if (dest!=0)  $fwrite(dest,"           TX CMD > $%h  =  (%d) - (%d) = (%b %b).\n",16'(cmd),8'(bh),8'(bl),8'(bh),8'(bl));
  @(negedge clk);
  TB_cmd_ena = 0;
  TB_cmd_in  = 16'(0);
WDT_COUNTER = WDT_RESET_TIME;
end
endtask
// ***********************************************************************************************************
// task script_set_xy(integer src, integer dest);
// Sets x&y[#] with values from script file.
// ***********************************************************************************************************
task script_set_xy(integer src, integer dest, integer ln);
begin
   integer r;
   string         xory,msg;
   logic          xory_bit;
   logic   [1:0]  pxy;
   logic   [11:0] xyd;
   logic   [15:0] cmd;

  while (WAIT_IDLE && (WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear

   r = $fscanf(src,"%s%d%d",xory,pxy,xyd);   // read command line parameters
   xory_bit = 0;
   if (xory=="Y" || xory=="y") xory_bit = 1; // Convert the X/Y string input into a bit.
   cmd = {1'b1,xory_bit,pxy,xyd};            // generate the CMD number

   $sformat(msg,"Set %s[%d] = %d.",(xory_bit ? "Y" : "X"),pxy,xyd); // Create the log and waveform message.
   //$sformat(msg,"Set %s[%d] = %d.",xory,pxy,xyd);                 // Create the log and waveform message.

   if (dest!=0) $fwrite(dest,"%s\n",msg);

   send_cmd(cmd,msg,ln,dest);
if (dest!=0) $fwrite(dest,"\n"); // Add a carrige return.
end
endtask

// ***********************************************************************************************************
// task set_xy(integer xory_bit,integer xyp, integer xyd);
// Sets x&y[#] with values from script file.
// ***********************************************************************************************************
task set_xy(logic xory_bit,logic unsigned [1:0] pxy, logic signed [11:0] xyd,string msg, integer line, integer dest);
begin
   logic   [15:0] cmd;
   cmd = {1'b1,xory_bit,pxy,xyd};  // generate the CMD number
   send_cmd(cmd,msg,line,dest);
end
endtask

// ***********************************************************************************************************
// task max_xy(integer src, integer dest);
// Sets maximum x&y drawing coordinates with values from script file.
// ***********************************************************************************************************
task max_xy(integer src, integer dest, integer ln);
begin
   integer r;
   string         msg;
   logic signed  [11:0] x,y;

  while (WAIT_IDLE && (WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear

   r = $fscanf(src,"%d%d",x,y);   // read command line parameters

   $sformat(msg,"Max(%d,%d).",x,y); // Create the log and waveform message.
   if (dest!=0) $fwrite(dest,"%s\n",msg);

   set_xy(0,3,x,msg,ln,dest);
   set_xy(1,3,y,msg,ln,dest);
   send_cmd({8'(92),8'(0)},msg,ln,dest);  // Command 93, copy XY[3] to max X/Y

//cmd_null( "" ); // Waits a clock & Leaves a clear space on the waveform
if (dest!=0) $fwrite(dest,"\n"); // Add a carrige return.

end
endtask


// ***********************************************************************************************************
// task set_paget(integer src, integer dest);
// Sets x&y[#] with values from script file.
// ***********************************************************************************************************
task set_paget(integer src, integer dest, integer ln);
begin

//logic unsigned [23:0] PAGER_base_adr[0:1]   = '{0,0}; // srce/dest base address.
//logic unsigned [23:0] PAGER_base_width[0:1] = '{0,0}; // srce/dest bitmap width.
//logic unsigned [ 7:0] PAGER_base_depth[0:1] = '{0,0}; // srce/dest bitmap depth.

   integer r;
   string         ssd,msg;
   logic          sd;
   logic   [15:0] cmd;

  while (WAIT_IDLE && (WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear

   r = $fscanf(src,"%s",ssd);                                                                // retrieve the SOURCE/DEST flag
   sd = 0;
   if (ssd[0]=="d" || ssd[0]=="D") sd = 1;                                                   // Convert the SOURCE/DEST string input into a bit.

   r = $fscanf(src,"%h%d%d",PAGER_base_adr[sd],PAGER_base_width[sd],PAGER_base_depth[sd]); // retrieve the SOURCE/DEST flag

   $sformat(msg,"SET_PAGET %s addr(h%h) width(%d) depth(%d)",(sd ? "Dest" : "Srce"),PAGER_base_adr[sd],16'(PAGER_base_width[sd]),5'(PAGER_base_depth[sd])); // Create the log and waveform message.

   if (dest!=0) $fwrite(dest,"%s\n",msg);


set_xy(1,2,PAGER_base_adr[sd][23:12]  ,msg, ln,dest);  // Store base address in XY[2]
set_xy(0,2,PAGER_base_adr[sd][11:0 ]  ,msg, ln,dest);
set_xy(1,3,PAGER_base_width[sd][23:12],msg, ln,dest);  // Store bitmap width in XY[3]
set_xy(0,3,PAGER_base_width[sd][11:0 ],msg, ln,dest);

send_cmd({5'b01111,1'(sd),2'(2),8'(PAGER_base_depth[sd]-1)},msg,ln,dest);  // Send set paget address using XY[2], includes bits/pixel depth
send_cmd({8'(112+sd),           8'(PAGER_base_depth[sd]-1)},msg,ln,dest);  // Send set paget width   using XY[3], includes bits/pixel depth

//cmd_null( "" ); // Waits a clock & Leaves a clear space on the waveform
if (dest!=0) $fwrite(dest,"\n"); // Add a carriage return.

end
endtask


// ***********************************************************************************************************
// task draw(integer src, integer dest, integer ln);
// Sets draw the selected shape
// ***********************************************************************************************************
task draw(integer src, integer dest, integer ln);
begin

   integer unsigned r,q1,q2;
   string         shape,msg;
   logic signed   [11:0] x [0:3];
   logic signed   [11:0] y [0:3];
   logic unsigned [7:0]  color ;
   logic                 fill;
   logic          [1:0]  quad;

   logic        [15:0] cmd;

  while (WAIT_IDLE && (WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear

   r = $fscanf(src,"%s",shape);                      // retrieve which shape to draw

case (shape[0]) // only analyze the first letter of the shape string.

   "p","P" : begin // draw a pixel
 
            r = $fscanf(src,"%d%d%d",x[0],y[0],color); // retrieve the SOURCE/DEST flag
            $sformat(msg,"Draw Pixel    (%d,%d), %d.",x[0],y[0],color); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);
             set_xy(0,0,x[0],msg,ln,dest);
             set_xy(1,0,y[0],msg,ln,dest);

             //        draw  fill  shape   color
             send_cmd({4'(0),1'(0),3'(1),8'(color)},msg,ln,dest);  // 1=draw pixel
             end

   "l","L" : begin // draw a line
 
            r = $fscanf(src,"%d%d%d%d%d",x[0],y[0],x[1],y[1],color); // retrieve the SOURCE/DEST flag
            $sformat(msg,"Draw Line     (%d,%d)-(%d,%d), %d.",x[0],y[0],x[1],y[1],color); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);
             set_xy(0,0,x[0],msg,ln,dest);
             set_xy(1,0,y[0],msg,ln,dest);
             set_xy(0,1,x[1],msg,ln,dest);
             set_xy(1,1,y[1],msg,ln,dest);

             //        draw  fill  shape   color
             send_cmd({4'(0),1'(0),3'(2),8'(color)},msg,ln,dest);  // 2=draw line
             end

   "b","B" : begin // draw a box
 
            r = $fscanf(src,"%d%d%d%d%d%d",x[0],y[0],x[1],y[1],color,fill); // retrieve the SOURCE/DEST flag
            $sformat(msg,"Draw Box      (%d,%d)-(%d,%d), %d%s",x[0],y[0],x[1],y[1],color,(fill ? ", filled. ":", no-fill.")); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);
             set_xy(0,0,x[0],msg,ln,dest);
             set_xy(1,0,y[0],msg,ln,dest);
             set_xy(0,1,x[1],msg,ln,dest);
             set_xy(1,1,y[1],msg,ln,dest);

             //        draw     fill  shape    color
             send_cmd({4'(0),1'(fill),3'(4),8'(color)},msg,ln,dest);  // 4=draw box
             end

   "t","T" : begin // draw a triangle
 
            r = $fscanf(src,"%d%d%d%d%d%d%d%d",x[0],y[0],x[1],y[1],x[2],y[2],color,fill); // retrieve the SOURCE/DEST flag
            $sformat(msg,"Draw Triangle (%d,%d)-(%d,%d)-(%d,%d), %d%s",x[0],y[0],x[1],y[1],x[2],y[2],color,(fill ? ", filled. ":", no-fill.")); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);
             set_xy(0,0,x[0],msg,ln,dest);
             set_xy(1,0,y[0],msg,ln,dest);
             set_xy(0,1,x[1],msg,ln,dest);
             set_xy(1,1,y[1],msg,ln,dest);
             set_xy(0,2,x[2],msg,ln,dest);
             set_xy(1,2,y[2],msg,ln,dest);

             //        draw     fill  shape    color
             send_cmd({4'(0),1'(fill),3'(3),8'(color)},msg,ln,dest);  // 3=draw triangle
             end

   "q","Q" : begin // draw a quadrilateral
 
            r = $fscanf(src,"%d%d%d%d%d%d%d%d%d%d",x[0],y[0],x[1],y[1],x[2],y[2],x[3],y[3],color,fill); // retrieve the SOURCE/DEST flag
            $sformat(msg,"Draw Quad     (%d,%d)-(%d,%d)-(%d,%d)-(%d,%d), %d%s",x[0],y[0],x[1],y[1],x[2],y[2],x[3],y[3],color,(fill ? ", filled. ":", no-fill.")); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);
             set_xy(0,0,x[0],msg,ln,dest);
             set_xy(1,0,y[0],msg,ln,dest);
             set_xy(0,1,x[1],msg,ln,dest);
             set_xy(1,1,y[1],msg,ln,dest);
             set_xy(0,2,x[2],msg,ln,dest);
             set_xy(1,2,y[2],msg,ln,dest);
             set_xy(0,3,x[3],msg,ln,dest);
             set_xy(1,3,y[3],msg,ln,dest);

             //        draw     fill  shape    color
// When filled, draw a filled triangle plus a filled quad, otherwise just draw a quad
if (fill)    send_cmd({4'(0),1'(fill),3'(3),8'(color)},msg,ln,dest);  // 3=draw triangle, *** When a quad is filled, you must send a filled triangle & a filled quad
             send_cmd({4'(0),1'(fill),3'(5),8'(color)},msg,ln,dest);  // 5=draw quad
             end


   "e","E" : begin // draw an Ellipse
 
            r = $fscanf(src,"%d%d%d%d%d%d%d",x[0],y[0],x[1],y[1],color,q2,fill); // retrieve the SOURCE/DEST flag
            $sformat(msg,"Draw Ellipse  P(%d,%d), R(%d,%d), C(%d), Q(%d), F(%d).",x[0],y[0],x[1],y[1],color,3'(q2),fill); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);
             set_xy(0,0,x[0],msg,ln,dest);
             set_xy(1,0,y[0],msg,ln,dest);
             set_xy(0,1,x[1],msg,ln,dest);
             set_xy(1,1,y[1],msg,ln,dest);

                 if (q2>3) begin    // setup for loop to draw all 4 quadrants
                           q1=0;
                           q2=4;
                 end else begin    // setup for loop to draw 1 quadrant
                           q1=q2;
                           q2=q2+1;
                 end

                 for (int unsigned q=q1 ; q<q2 ; q++ ) begin // setup loop to draw the requested quadrants.

                 while (WAIT_IDLE && (WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear
                $sformat(msg,"Draw Ellipse  C(%d,%d), R(%d,%d), C(%d), Q(%d), F(%d).",x[0],y[0],x[1],y[1],color,3'(q),fill); // Create the log and waveform message.
                 send_cmd({8'(7)               ,6'(0),2'(q)},msg,ln,dest); // 7 = (lower 2 bits) = select ellipse quadrant.
                 send_cmd({4'(0),1'(fill),3'(6),8'(color)  },msg,ln,dest);   // 6 = draw ellipse

                 end
             end

   default : begin
                 while ((WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear
                  $sformat(msg,"Unknown draw shape '%s' at line number %d.\nProcessign stopped due to error.\n",shape,13'(ln));
                  $display("%s",msg);
                  cmd_null( msg ); // Waits a clock & Leaves a clear space on the waveform
                  while ((WDT_COUNTER >= 2 )) @(negedge clk); // wait for busy to clear
                  if (dest!=0) $fwrite(dest,"%s",msg);
                  $stop;

             end


endcase

//cmd_null( "" ); // Waits a clock & Leaves a clear space on the waveform
if (dest!=0) $fwrite(dest,"\n"); // Add a carriage return.

end
endtask


// ***********************************************************************************************************
// task load_gpu_ram(integer src,dest,line_number,endian);
// Sets draw the selected shape
// ***********************************************************************************************************

task load_gpu_ram(integer src,dest,line_number,endian);
begin

    string                  bin_file_name, msg;
    integer unsigned        bin_src, mem_adr, max_adr, r;
    logic unsigned [7:0]    byte_h,byte_l;

    max_adr = (2**(PIXIE_MEM_ADR-1));

    wait_idle();

    r = $fscanf(src,"%s",bin_file_name);                      // retrieve which shape to draw

    bin_src = $fopen(bin_file_name,"rb");
    if (bin_src==0)
    begin
       $display("Could not open file '%s' for reading.",bin_file_name);
       $stop;     
    end
    $display(" *************************************************************** ");
    $display(" *** LOAD_GPU_RAM '%s' into GPU RAM. ***** ",bin_file_name);
    $display(" *************************************************************** ");

                 $sformat(msg,"LOAD_GPU_RAM %s.",bin_file_name);
                 cmd_null(msg);
                 cmd_null(msg);
                 if (dest!=0) $fwrite(dest,"%s\n",msg);


for (mem_adr = 0 ; ((mem_adr < max_adr) && (! $feof(bin_src))) ; mem_adr ++ ) begin
          byte_h = $fgetc(bin_src);
          byte_l = $fgetc(bin_src);
          if (! $feof(bin_src)) begin
               if (endian == 0) GPU_RAM[mem_adr] = {byte_h,byte_l};
               else             GPU_RAM[mem_adr] = {byte_l,byte_h};
          end
          end

    $fclose(bin_src);
end
endtask

// ***********************************************************************************************************
// task load_gpu_ram(integer src,dest,line_number,endian);
// Sets draw the selected shape
// ***********************************************************************************************************

task save_gpu_ram(integer src,dest,line_number,endian);
begin

    string                  bin_file_name, msg;
    integer unsigned        bin_src, mem_adr, max_adr, r;
    logic unsigned [7:0]    b [3:0];

    max_adr = (2**(PIXIE_MEM_ADR-1));

    wait_idle();

    r = $fscanf(src,"%s",bin_file_name);                      // retrieve which shape to draw

    bin_src = $fopen(bin_file_name,"wb");
    if (bin_src==0)
    begin
       $display("Could not open file '%s' for writing.",bin_file_name);
       $stop;     
    end
    $display(" *************************************************************** ");
    $display(" *** SAVE_GPU_RAM to file '%s'. ***** ",bin_file_name);
    $display(" *************************************************************** ");

                 $sformat(msg,"SAVE_GPU_RAM %s.",bin_file_name);
                 cmd_null(msg);
                 cmd_null(msg);
                 if (dest!=0) $fwrite(dest,"%s\n",msg);


     for (mem_adr = 0 ; mem_adr < max_adr ; mem_adr +=2 ) begin

          b[0] = GPU_RAM[mem_adr+0][15:8];
          b[1] = GPU_RAM[mem_adr+0][7:0];
          b[2] = GPU_RAM[mem_adr+1][15:8];
          b[3] = GPU_RAM[mem_adr+1][7:0];

          if (endian == 0) $fwrite(bin_src,"%u",{b[3],b[2],b[1],b[0]});
          else             $fwrite(bin_src,"%u",{b[0],b[1],b[2],b[3]});

     end

    $fclose(bin_src);
end
endtask


// ***********************************************************************************************************
// function logic unsigned [7:0] pixie_pixel (bit z,logic unsigned [11:0] x,y);
// Reads GPU memory and returns a PIXEL, basically emulates MAGGIE/BART, or core of PIXIE
// ***********************************************************************************************************

function logic unsigned [7:0] pixie_pixel (bit z,logic unsigned [11:0] x,y);

logic [2:0]  LUT_bits_to_shift[0:15] ;  // shift bits/pixel-1  0=1 bit, 1=2bit, 3=4bit, 7=8bit, 15-16bit.
logic [3:0]  LUT_shift [0:255]       ;
logic [15:0] LUT_mask  [0:15]        ;  // mask result bits after shift pixel-1  0=1 bit, 1=2bit, 3=4bit, 7=8bit, 15-16bit.

logic unsigned [7:0] color_gain [0:15] ;     // Amplifies the color number of lower bitplane displays
logic unsigned [(PIXIE_MEM_ADR-1):0] raddr;
logic unsigned [3:0] sb ;


LUT_shift = '{
15,14,13,12,11,10, 9, 8, 7, 6, 5, 4, 3, 2, 1, 0,  // Shift values for bpp=0, target=0 through 15.
14,12,10, 8, 6, 4, 2, 0,14,12,10, 8, 6, 4, 2, 0,  // Shift values for bpp=1, target=0 through 15.
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=2, invalid bitplane mode, no shift
12, 8, 4, 0,12, 8, 4, 0,12, 8, 4, 0,12, 8, 4, 0,  // Shift values for bpp=3, target=0 through 15.
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=4, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=5, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=6, invalid bitplane mode, no shift
 8, 0, 8, 0, 8, 0, 8, 0, 8, 0, 8, 0, 8, 0, 8, 0,  // Shift values for bpp=7, target=0 through 15.
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=8, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=9, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=10, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=11, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=12, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=13, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,  // Shift values for bpp=14, invalid bitplane mode, no shift
 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0   // Shift values for bpp=15, target=0 through 15.
};

LUT_bits_to_shift  = '{  4,  3,  3,  2,  2,  2,  2,  1,  1,  1,  1,  1,  1,  1,  1,    0 }; // shift bits/pixel-1  0=1 bit, 1=2bit, 3=4bit, 7=8bit, 15-16bit.
LUT_mask           = '{  1,  3,  3, 15, 15, 15, 15,255,255,255,255,255,255,255,255,65535 }; // mask result bits after shift pixel-1  0=1 bit, 1=2bit, 3=4bit, 7=8bit, 15-16bit.
color_gain         = '{255, 63, 63, 15, 15, 15, 15,  1,  1,  1,  1,  1,  1,  1,  1,    1 }; // Amplifies the color number of lower bitplane displays

    sb    =  PAGER_base_depth[z] - 1 ;
    raddr =  PAGER_base_adr[z]   + (y * PAGER_base_width[z]) + x ; // calculate the read address.

    return 8'(  (( GPU_RAM[raddr >> LUT_bits_to_shift[sb]] >> LUT_shift[{sb,raddr[3:0]}] )  & LUT_mask[sb]  )   * color_gain[sb] );

endfunction




// ***********************************************************************************************************
// task draw(integer src, integer dest, integer ln);
// Sets draw the selected shape
// ***********************************************************************************************************
task blit(integer src, integer dest, integer ln);
begin

   integer unsigned r,q1,q2;
   string         func,msg;
   logic unsigned [11:0] x [0:3];
   logic unsigned [11:0] y [0:3];
   logic unsigned [7:0]  color ;
   logic                 fill;
   logic          [1:0]  quad;

   real           usx,usy,dsx,dsy;

   logic          [15:0] cmd;

  while (WAIT_IDLE && (WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear

   r = $fscanf(src,"%s",func);                      // retrieve which shape to draw

case (func[0]) // only analyze the first letter of the shape string.

   "c","C" : begin // Set blitter config.
 
            r = $fscanf(src,"%b%b%b%b%b%b%b%b",color[0],color[1],color[2],color[3],color[4],color[5],color[6],color[7]);       // retrieve transparent color
            $sformat(msg,"BLIT config ena %b,msk %b,hc %b,mir %b,vc %b,flp %b,r90 %b,r45 %b.",color[0],color[1],color[2],color[3],color[4],color[5],color[6],color[7]); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);

             //        draw   func    color
             send_cmd({4'(0),4'(0),8'(color)},msg,ln,dest);  // 0=set the blitter transparency mask color
             end

   "t","T" : begin // Select transparent color.
 
            r = $fscanf(src,"%d",color);                           // retrieve transparent color
            $sformat(msg,"BLIT t-color %d.",color); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);

             //        draw   func    color
             send_cmd({4'(0),4'(8),8'(color)},msg,ln,dest);  // 8=set the blitter transparency mask color
             end

   "p","P" : begin // set source image position and size
 
            r = $fscanf(src,"%d%d%d%d",x[2],y[2],x[3],y[3]);                           // retrieve transparent color
            $sformat(msg,"BLIT source pos(%d,%d), size(%d,%d).",x[2],y[2],x[3],y[3]); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);

            //x[3]=x[3]-1; // *** Width and height need to be subtracted by 1.
            //y[3]=y[3]-1;

             set_xy(0,2,x[2],msg,ln,dest);
             set_xy(1,2,y[2],msg,ln,dest);
             set_xy(0,3,x[3],msg,ln,dest);
             set_xy(1,3,y[3],msg,ln,dest);


             //         func    N/A
             send_cmd({8'(118),8'(0)},msg,ln,dest);  // 118 = transfer xy[2] to blitter source offset X&Y position
             send_cmd({8'(117),8'(0)},msg,ln,dest);  // 117 = transfer xy[3] to blitter copy width and height
             end


   "s","S" : begin // Sets the blitter scale.
 
            r = $fscanf(src,"%f%f%f%f",usx,usy,dsx,dsy);                           // retrieve transparent color

            if (usx>4095.0)   usx  = 4095.0;         // cap and limit input us-sample scale
                              x[0] = int'(4096/usx);
            if (usx<=1.0)     x[0] = 0;              // 1.00000 is a special case where us(X/Y) =0
            if (usx<=1.0)     usx  = 1.0;
            if (usy>4095.0)   usy  = 4095.0;         // cap and limit input us-sample scale
                              y[0] = int'(4096/usy);
            if (usy<=1.0)     y[0] = 0;              // 1.00000 is a special case where us(X/Y) =0
            if (usy<=1.0)     usy  = 1.0;

            if (dsx<0.000245) dsx  = 0.000245;       // cap and limit input down-sample scale
                              x[1] = int'(4096*dsx);
            if (dsx>=1.0)     x[1] = 0;              // 1.00000 is a special case where ds(X/Y) =0
            if (dsx>=1.0)     dsx  = 1.0;
            if (dsy<0.000245) dsy  = 0.000245;       // cap and limit input down-sample scale
                              y[1] = int'(4096*dsy);
            if (dsy>=1.0)     y[1] = 0;              // 1.00000 is a special case where ds(X/Y) =0
            if (dsy>=1.0)     dsy  = 1.0;


            $sformat(msg,"BLIT SCALE us(%f,%f), ds(%f,%f).",usx,usy,dsx,dsy); // Create the log and waveform message.

            if (dest!=0) $fwrite(dest,"%s UpSamp=(%d,%d)/4096, DownSamp=(%d,%d)/4096. *(0=4096).\n",msg,x[0],y[0],x[1],y[1]);

             set_xy(0,0,x[0],msg,ln,dest);
             set_xy(1,0,y[0],msg,ln,dest);
             set_xy(0,1,x[1],msg,ln,dest);
             set_xy(1,1,y[1],msg,ln,dest);

             //         Draw  Set Blit Scale
             send_cmd({8'(9),8'(3)},msg,ln,dest);  // 9 = Draw func set blit scale, 3 = set src&dest scale with xy[0],xy[1]
             end


   default : begin
                 while ((WDT_COUNTER > SYS_IDLE_TIME)) @(negedge clk); // wait for busy to clear
                  $sformat(msg,"Unknown BLIT function '%s' at line number %d.\nProcessign stopped due to error.\n",func,13'(ln));
                  $display("%s",msg);
                  cmd_null( msg ); // Waits a clock & Leaves a clear space on the waveform
                  while ((WDT_COUNTER >= 2 )) @(negedge clk); // wait for busy to clear
                  if (dest!=0) $fwrite(dest,"%s",msg);
                  $stop;

             end


endcase

//cmd_null( "" ); // Waits a clock & Leaves a clear space on the waveform
if (dest!=0) $fwrite(dest,"\n"); // Add a carriage return.

end
endtask

// ***********************************************************************************************************
// task vwait(integer src, integer dest, integer ln);
// Sets the VWAIT routine.
// ***********************************************************************************************************
task vwait(integer src, integer dest, integer ln);
begin

   integer unsigned        r;
   string                  msg;
   logic   unsigned [3:0]  framew ;
   logic   unsigned [7:0]  linew ;
   logic   unsigned [7:0]  cmd;

 
            r = $fscanf(src,"%d%d",framew,linew);       // retrieve number of frames to wait & which video line to wait for.

            $sformat(msg,"VWAIT for %d frames, until line number %d.",framew,linew); // Create the log and waveform message.
            if (dest!=0) $fwrite(dest,"%s\n",msg);


             send_cmd({8'(15),8'(linew)},msg,ln,dest);  // Which video line to wait for.
             cmd = 8'b10000000 | framew;                // Set the frame count and multiply the video line to wait for by 1.
             send_cmd({8'( 7),8'(cmd  )},msg,ln,dest);  // Send the wait command with frame count.

end
endtask

endmodule
